`ifndef WISHBONE_DEFS_SVH
`define WISHBONE_DEFS_SVH

typedef enum logic {
    IDLE,
    BUS_WAIT
} master_state_t;

`endif
